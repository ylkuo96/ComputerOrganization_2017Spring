module opUnit(
    output wire result,
    output wire carryout,
    input wire [31:0]a,b,
    input wire carryin,
    input wire less, 
);

endmodule
