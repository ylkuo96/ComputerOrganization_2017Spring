module alu(
    output [31:0]result, 
    output [31:0] result,
    output zero,
    output cout,

    input rst_n,
    input [31:0] a, b,
    input [3:0] ALU_control,
);
/*
output wire result,
    output wire carryout,
    input wire [31: 0]a,b,
    input wire [3:0] opcode,
    input wire carryin,
    input wire less, 
*/


opUnit u1( );


endmodule
